// Computer Architecture (CO224) - Lab 05
// Design: Testbench of Integrated CPU of Simple Processor
// Author: Isuru Nawinne
`include "cpu.v"
`include "imemory.v"
`include "icache.v"
`timescale 1ns/1ps
module cpu_tb;

    reg CLK, RESET;
    wire [31:0] PC;
    wire [31:0] INSTRUCTION;
    wire BUSYWAIT;

    /* 
    ------------------------
     SIMPLE INSTRUCTION MEM
    ------------------------
    */
    
    // TODO: Initialize an array of registers (8x1024) named 'instr_mem' to be used as instruction memory
    
    // TODO: Create combinational logic to support CPU instruction fetching, given the Program Counter(PC) value 
    //       (make sure you include the delay for instruction fetching here)
    reg [7:0] instr_mem[1023:0];
     //assign #2 INSTRUCTION={instr_mem[PC+3], instr_mem[PC+2], instr_mem[PC+1], instr_mem[PC]};
    initial
    begin
        // Initialize instruction memory with the set of instructions you need execute on CPU
        
        // METHOD 1: manually loading instructions to instr_mem
        // {instr_mem[10'd3], instr_mem[10'd2], instr_mem[10'd1], instr_mem[10'd0]} = 32'b00000000000001000000000000000101;
        // {instr_mem[10'd7], instr_mem[10'd6], instr_mem[10'd5], instr_mem[10'd4]} = 32'b00000000000000100000000000001001;
        // {instr_mem[10'd11], instr_mem[10'd10], instr_mem[10'd9], instr_mem[10'd8]} = 32'b00000010000001100000010000000010;
        
        // METHOD 2: loading instr_mem content from instr_mem.mem file
        $readmemb("instr_mem.mem", instr_mem);
    end
    
    
    
    /* 
    -----
     CPU
    -----
    */
    wire MEM_BUSYWAIT,MEME_READ;
    wire [127:0]MEM_INSTRUCTION;
    wire [5:0]MEM_ADDRESS;
    icache myicache(BUSYWAIT,CLK,RESET, INSTRUCTION, PC[9:2],MEM_BUSYWAIT,MEM_INSTRUCTION,MEM_READ,MEM_ADDRESS);
    instruction_memory myimem(CLK,MEM_READ,MEM_ADDRESS,MEM_INSTRUCTION,MEM_BUSYWAIT);
    cpu mycpu( INSTRUCTION, CLK, RESET,PC,BUSYWAIT);
    integer i;
    initial
    begin
    
        // generate files needed to plot the waveform using GTKWave
        $dumpfile("cpu_wavedata.vcd");
		$dumpvars(0, cpu_tb);
        
        for (i=0 ;i<8;i=i+1)
            $dumpvars(1,cpu_tb.mycpu.reg_8x8.regArr[i]);
        for(i=0;i<256;i++)
            $dumpvars(1,cpu_tb.mycpu.dm2.memory_array[i]);
        for(i=0;i<8;i++)
            $dumpvars(1,cpu_tb.mycpu.dcache_cpu.cache_array[i]);
        for(i=0;i<8;i++)
            $dumpvars(1,cpu_tb.myicache.icache_array[i]);
        for(i=0;i<1024;i++)
            $dumpvars(1,cpu_tb.myimem.memory_array[i]);
        for(i=0;i<8;i++)
            $dumpvars(1,cpu_tb.myicache.valid_array[i]);
        for(i=0;i<8;i++)
            $dumpvars(1,cpu_tb.myicache.tag_array[i]);
        CLK = 1'b0;
        RESET = 1'b0;
        
        // TODO: Reset the CPU (by giving a pulse to RESET signal) to start the program execution
        RESET = 1'b1;
        #6
        RESET = 1'b0;
        // finish simulation after some time
        #2900
        $finish;
        
    end
    
    // clock signal generation
    always
        #4 CLK = ~CLK;
        

endmodule